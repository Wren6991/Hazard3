// Minimal Hazard3 config for testbench

localparam RESET_VECTOR        = 32'h40;
localparam MTVEC_INIT          = 32'h0;
localparam EXTENSION_A         = 0;
localparam EXTENSION_C         = 0;
localparam EXTENSION_M         = 0;
localparam EXTENSION_ZBA       = 0;
localparam EXTENSION_ZBB       = 0;
localparam EXTENSION_ZBC       = 0;
localparam EXTENSION_ZBS       = 0;
localparam EXTENSION_ZBKB      = 0;
localparam EXTENSION_ZIFENCEI  = 0;
localparam EXTENSION_XH3BEXTM  = 0;
localparam EXTENSION_XH3IRQ    = 0;
localparam EXTENSION_XH3PMPM   = 0;
localparam EXTENSION_XH3POWER  = 0;
localparam CSR_M_MANDATORY     = 1;
localparam CSR_M_TRAP          = 1;
localparam CSR_COUNTER         = 0;
localparam U_MODE              = 0;
localparam PMP_REGIONS         = 0;
localparam PMP_GRAIN           = 0;
localparam PMP_HARDWIRED       = {PMP_REGIONS{1'b0}};
localparam PMP_HARDWIRED_ADDR  = {PMP_REGIONS{32'h0}};
localparam PMP_HARDWIRED_CFG   = {PMP_REGIONS{8'h00}};
localparam DEBUG_SUPPORT       = 0;
localparam BREAKPOINT_TRIGGERS = 4;
localparam NUM_IRQS            = 32;
localparam IRQ_PRIORITY_BITS   = 0;
localparam IRQ_INPUT_BYPASS    = {NUM_IRQS{1'b0}};
localparam MVENDORID_VAL       = 32'hdeadbeef;
localparam MIMPID_VAL          = 32'h12345678;
localparam MHARTID_VAL         = 32'h9abcdef0;
localparam MCONFIGPTR_VAL      = 32'h0;
localparam REDUCED_BYPASS      = 1;
localparam MULDIV_UNROLL       = 1;
localparam MUL_FAST            = 0;
localparam MUL_FASTER          = 0;
localparam MULH_FAST           = 0;
localparam FAST_BRANCHCMP      = 0;
localparam RESET_REGFILE       = 1;
localparam BRANCH_PREDICTOR    = 0;
localparam MTVEC_WMASK         = 32'hfffffffd;
